//-------------------------------------------------------------------------------------------------
//  File name	  	: aes_mixcolumn.v
//  Project		: AES128
//  Author		: Do Quang Huy
//  Description		: Round Contants 
//
//  Referents		: Pham Hoai Luan.
//-------------------------------------------------------------------------------------------------


module aes_inv_mixcolumn(
	inv_mixcolumn_in,
	inv_mixcolumn_out
);

//---------------------------------------------------------------------------------------------
//  Ports
//---------------------------------------------------------------------------------------------

  input  wire [31:0] inv_mixcolumn_in;
  output wire [31:0] inv_mixcolumn_out;
  
//----------------------------------------------------------------
// Architecture:  Controlling the value output
//----------------------------------------------------------------
  assign inv_mixcolumn_out = inv_mixw(inv_mixcolumn_in);
  
//----------------------------------------------------------------
//  Architecture:  Controlling the value output
//----------------------------------------------------------------

// This operation on bytes is denoted by gm().
// Multiplication by higher powers of x can be implemented by repeated application of gm().
// By adding intermediate results, multiplication by any constant can be implemented. 
// {57} ? {02} = gm({57}) = {ae}
// {57} ? {04} = gm({ae}) = {47}
// {57} ? {08} = gm({47}) = {8e}
// {57} ? {10} = gm({8e}) = {07}
// {57} ? {13} = {57} ? ({01} ^ {02} ^ {10})
// = {57} ^ {ae} ^ {07}
// = {fe}.  

function [7 : 0] gm2(input [7 : 0] op);
    begin
      gm2 = {op[6 : 0], 1'b0} ^ (8'h1b & {8{op[7]}});
    end
  endfunction // gm2

  function [7 : 0] gm3(input [7 : 0] op);
    begin
      gm3 = gm2(op) ^ op;
    end
  endfunction // gm3

  function [7 : 0] gm4(input [7 : 0] op);
    begin
      gm4 = gm2(gm2(op));
    end
  endfunction // gm4

  function [7 : 0] gm8(input [7 : 0] op);
    begin
      gm8 = gm2(gm4(op));
    end
  endfunction // gm8

  function [7 : 0] gm09(input [7 : 0] op);
    begin
      gm09 = gm8(op) ^ op;
    end
  endfunction // gm09

  function [7 : 0] gm11(input [7 : 0] op);
    begin
      gm11 = gm8(op) ^ gm2(op) ^ op;
    end
  endfunction // gm11

  function [7 : 0] gm13(input [7 : 0] op);
    begin
      gm13 = gm8(op) ^ gm4(op) ^ op;
    end
  endfunction // gm13

  function [7 : 0] gm14(input [7 : 0] op);
    begin
      gm14 = gm8(op) ^ gm4(op) ^ gm2(op);
    end
  endfunction // gm14

  function [31 : 0] inv_mixw(input [31 : 0] w);
    reg [7 : 0] b0, b1, b2, b3;
    reg [7 : 0] mb0, mb1, mb2, mb3;
    begin
      b0 = w[31 : 24];
      b1 = w[23 : 16];
      b2 = w[15 : 08];
      b3 = w[07 : 00];

      mb0 = gm14(b0) ^ gm11(b1) ^ gm13(b2) ^ gm09(b3);
      mb1 = gm09(b0) ^ gm14(b1) ^ gm11(b2) ^ gm13(b3);
      mb2 = gm13(b0) ^ gm09(b1) ^ gm14(b2) ^ gm11(b3);
      mb3 = gm11(b0) ^ gm13(b1) ^ gm09(b2) ^ gm14(b3);

      inv_mixw = {mb0, mb1, mb2, mb3};
    end
  endfunction
endmodule 


